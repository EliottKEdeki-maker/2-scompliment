`timescale 1ns / 1ps
module invert();

  input
  output
  wire
