`timescale 1ns / 1ps
module invert(x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11;);

  input x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,d,j,k,t_clk;
  output q1,q2;
  wire dp1,s,r,dp2, jk1, jk2, jk3;

  
