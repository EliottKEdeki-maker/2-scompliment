`timescale 1ns / 1ps
module invert(x,r,q1,q2);

  input x1,x2,x3,r;
  output q1, q2, o1;
  wire
