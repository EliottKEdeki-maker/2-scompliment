`timescale 1ns / 1ps
module invert();

  input x,r;
  output q1, q2;
  wire
