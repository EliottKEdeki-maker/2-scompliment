`timescale 1ns / 1ps
module invert(x,r,q1,q2);

  input x,r;
  output q1, q2;
  wire
